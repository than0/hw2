package global_types;
//define the rounding modes used by the modules
typedef enum logic [2:0] {IEEE_near, IEEE_zero, IEEE_pinf, IEEE_ninf, near_up, away_zero} rounding_mode;

//define the random edge cases for testing
typedef enum logic [31:0] {pos_qnan = 32'b01111111101100100100001001110111, neg_qnan = 32'b11111111101000111011001000110110,
				pos_snan = 32'b01111111110011010001101011101100, neg_snan = 32'b11111111110100001010011101010001,
				pos_inf = 32'b01111111100000000000000000000000, neg_inf = 32'b11111111100000000000000000000000,
				pos_zero = 32'b00000000000000000000000000000000, neg_zero = 32'b10000000000000000000000000000000,
			        pos_denorm = 32'b00000000001011011010010110110010, neg_denorm = 32'b10000000010100001110110111001101,
				pos_norm = 32'b01001101110100010101111001001101, neg_norm = 32'b11001110101100101101100101011001} boundary_cond;

endpackage
